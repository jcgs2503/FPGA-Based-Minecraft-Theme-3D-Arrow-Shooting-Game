module texture_1_palette (
	input logic [7:0] index,
	output logic [3:0] red, green, blue
);

localparam [0:255][11:0] palette = {
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hD, 4'hD, 4'hC},
	{4'hD, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hD, 4'hD, 4'hC},
	{4'hD, 4'hD, 4'hC},
	{4'hD, 4'hD, 4'hC},
	{4'hD, 4'hD, 4'hC},
	{4'hD, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hE, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hD, 4'hD, 4'hC},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD},
	{4'hE, 4'hD, 4'hD}
};

assign {red, green, blue} = palette[index];

endmodule
